module input_output(input in, output out);
  assign out=1'b1;
  //assign out=in;
endmodule
